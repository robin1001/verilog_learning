module hello_world ();
    initial begin
        $display("hello world");
        $finish;
    end
endmodule
